Library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
entity DIEUKHIEN_CHOPHEP is
	Port ( CKHT,RST: in STD_LOGIC;
			 ENA_DB_1, ENA_DB_2: IN STD_LOGIC;
				OE: out STD_LOGIC_VECTOR (1 downto 0));
end DIEUKHIEN_CHOPHEP;
architecture Behavioral of DIEUKHIEN_CHOPHEP is
SIGNAL DEM_REG, DEM_NEXT: INTEGER RANGE 0 TO 9999:=0;
SIGNAL ENA_DB: STD_LOGIC;
begin
	PROCESS(CKHT,RST)
	BEGIN
	-- REGISTER FF-D
		IF (RST ='1') THEN DEM_REG <= 0;
		ELSIF FALLING_EDGE(CKHT) THEN DEM_REG <= DEM_NEXT;
		END IF;
	END PROCESS;
	-- DEM DEN LAN 31 THI RESET NEU KO THI DEM TIEP
	DEM_NEXT <= DEM_REG WHEN DEM_REG = 80 AND ENA_DB = '1' ELSE
	DEM_REG + 1 WHEN ENA_DB = '1' ELSE
	DEM_REG;
	PROCESS(DEM_REG, RST)
	BEGIN
		OE <= "00";
		IF RST = '1' THEN OE <= "00";
		ELSIF DEM_REG < 60 THEN OE <= "01";ENA_DB <= ENA_DB_1;
		ELSIF DEM_REG < 80 THEN OE <= "10";ENA_DB <= ENA_DB_2;
		END IF;
	END PROCESS;
end Behavioral;