-- CHUONG TRINH CON DA HOP 4 KENH 1 BIT

