
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity LED_STD_PST is
    Port (CKHT, RST, OE, ENA_DB:   in      STD_LOGIC;
				SO_LED :IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    		Q:      out     STD_LOGIC_VECTOR (7 downto 0));
end LED_STD_PST;

architecture Behavioral of LED_STD_PST is
SIGNAL 	Q_REG, Q_NEXT,X: STD_LOGIC_VECTOR(7 DOWNTO 0);
Begin
   PROCESS (CKHT, RST)
   BEGIN   
		IF  RST='1'             THEN    Q_REG	<=	(OTHERS => '0'); 
      ELSIF   FALLING_EDGE (CKHT)   THEN    Q_REG	<=	Q_NEXT;	
		END IF;
	END PROCESS;
X<= Q_REG(6 DOWNTO 0) & NOT Q_REG(7 )  WHEN SO_LED ="0001" 		  ELSE
	"00000000" WHEN SO_LED ="0011" AND Q_REG ="10000000"			  ELSE
	"11111111" WHEN SO_LED ="0011" AND Q_REG ="01111111" 			  ELSE 
	Q_REG(5 DOWNTO 0) & NOT Q_REG(7 DOWNTO 6) WHEN SO_LED ="0011" ELSE
	"00000000" WHEN SO_LED ="0111" AND (Q_REG ="11000000"OR Q_REG = "10000000") 	ELSE
	"11111111" WHEN SO_LED ="0111" AND (Q_REG ="01111111"OR Q_REG ="00111111") 	ELSE
	Q_REG(4 DOWNTO 0) & NOT Q_REG(7 DOWNTO 5 ) WHEN SO_LED ="0111" 					ELSE
	"00000000" WHEN SO_LED ="1111" AND (Q_REG ="11000000"OR Q_REG="10000000"OR  Q_REG= "11100000") 	ELSE
	"11111111" WHEN SO_LED ="1111" AND (Q_REG ="01111111"OR Q_REG ="00111111"OR Q_REG ="00011111")  ELSE
	Q_REG(3 DOWNTO 0) & NOT Q_REG(7 DOWNTO 4) ;
	
Q_NEXT  <=  (OTHERS => '0')			WHEN OE = '0' 		ELSE
				    X 						WHEN ENA_DB = '1' ELSE	
					Q_REG;					
Q <= Q_REG 									WHEN OE = '1' ELSE 
	(OTHERS => '0'); 
      
end Behavioral;

