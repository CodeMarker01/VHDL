library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity DK_8LED_2CT_AU_SANGDON is
	Port ( CKHT, BTN_N0: in STD_LOGIC;
			LED: out STD_LOGIC_VECTOR (7 downto 0));
end DK_8LED_2CT_AU_SANGDON;

architecture Behavioral of DK_8LED_2CT_AU_SANGDON is
SIGNAL ENA_DB, RST: STD_LOGIC;
SIGNAL Q_SD_PST, Q_SD_TSP: STD_LOGIC_VECTOR (7 downto 0);
SIGNAL OE: STD_LOGIC_VECTOR(1 DOWNTO 0);
Begin
	RST <= NOT BTN_N0;
CHIA_10ENA: ENTITY WORK.CHIA_10ENA
	PORT MAP ( CKHT => CKHT,
	ENA5HZ => ENA_DB);
LED_SANGDON_PST: ENTITY WORK.LED_SANGDON_PST
	PORT MAP ( CKHT => CKHT,
	RST => RST,
	ENA_DB => ENA_DB,
	OE => OE(0),
	Q => Q_SD_PST);
LED_SANGDON_TSP: ENTITY WORK.LED_SANGDON_TSP
	PORT MAP ( CKHT => CKHT,
	RST => RST,
	ENA_DB => ENA_DB,
	OE => OE(1),
	Q => Q_SD_TSP);
	DIEUKHIEN_CHOPHEP: ENTITY WORK.DIEUKHIEN_CHOPHEP
	PORT MAP ( CKHT => CKHT,
	RST => RST,
	ENA_DB => ENA_DB,
	OE => OE);
	
	LED <= Q_SD_TSP OR Q_SD_PST;
end Behavioral;