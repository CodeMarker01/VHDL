LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY DEM_8BIT IS
	PORT(CKHT,RST, BTN1,BTN2,BTN3,ENA1HZ,ENA5HZ:IN STD_LOGIC;			
			ENA_DB,HUONG,LED_HUONG,LED_XUNG,SS: OUT STD_LOGIC		
			);
END DEM_8BIT;

ARCHITECTURE BEHAVIORAL OF DEM_8BIT IS
SIGNAL Q1_REG,Q1_NEXT : STD_LOGIC;
SIGNAL Q2_REG,Q2_NEXT : STD_LOGIC;
SIGNAL Q3_REG,Q3_NEXT : STD_LOGIC;
BEGIN
	PROCESS(CKHT,RST)
	BEGIN
		IF RST='1' THEN Q1_REG <= '0';
							 Q2_REG <= '0';
							 Q3_REG <= '0';
		ELSIF FALLING_EDGE(CKHT) THEN 
											Q1_REG <= Q1_NEXT;
											Q2_REG <= Q2_NEXT;
											Q3_REG <= Q3_NEXT;
		END IF;
	END PROCESS;
	Q1_NEXT <=   	NOT Q1_REG	WHEN BTN1='1' ELSE
			         Q1_REG;	
	Q2_NEXT <=   	NOT Q2_REG		WHEN BTN2='1' ELSE
			         Q2_REG;
	Q3_NEXT <=   	NOT Q3_REG		WHEN BTN3='1' ELSE
			         Q3_REG;	
	ENA_DB 		<= ENA1HZ 	WHEN Q1_REG='0' ELSE ENA5HZ	;
	LED_XUNG		<=	'0' 		WHEN Q1_REG='0' ELSE '1'	;
	HUONG 		<= '0' 		WHEN Q2_REG='0' ELSE '1'	;	
	SS		 		<= '0' 	  	WHEN Q3_REG='0' ELSE '1';			
	LED_HUONG	<= '0' 		WHEN Q2_REG='0' ELSE '1'	;
	
	
END BEHAVIORAL;