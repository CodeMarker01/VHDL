
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;


entity XULY_MOD_DAUCHAM_NHAP_NHAY is
    Port ( CKHT, ENA_DB, ENA2HZ, ENA_UP, ENA_DW, ENA_NN, ENA_SS : in  STD_LOGIC;
           GIATRI_MOD : in  STD_LOGIC_VECTOR (1 downto 0);
           ENA_GIAIMA_8LED : out  STD_LOGIC_VECTOR (7 downto 0);
           DAU_CHAM_8LED : out  STD_LOGIC_VECTOR (7 downto 0));
end XULY_MOD_DAUCHAM_NHAP_NHAY;

architecture Behavioral of XULY_MOD_DAUCHAM_NHAP_NHAY is

SIGNAL ENAGM_8LED_REG: STD_LOGIC_VECTOR( 7 DOWNTO 0):=X"FF";
SIGNAL ENAGM_8LED_NEXT: STD_LOGIC_VECTOR( 7 DOWNTO 0);


begin
	PROCESS(CKHT)
	BEGIN
		IF FALLING_EDGE(CKHT) THEN 
											ENAGM_8LED_REG <= ENAGM_8LED_NEXT;
											
		END IF;
	END PROCESS;
	
	PROCESS(GIATRI_MOD, ENA2HZ, ENAGM_8LED_REG)
	BEGIN
		ENAGM_8LED_NEXT <= ENAGM_8LED_REG;
			IF (ENA_NN= '0' AND ENA_SS = '1' ) THEN
				IF ENA2HZ = '1' THEN 
					ENAGM_8LED_NEXT <= "000" & NOT ENAGM_8LED_REG( 4 DOWNTO 3) & '0' & NOT ENAGM_8LED_REG( 1 DOWNTO 0); --NHAP NHAY 2 LED GIAY
				END IF;
		ELSE 
			ENAGM_8LED_NEXT <= "00011011";
		END IF;
		END PROCESS;
		
		------------------------------------------------------------
	PROCESS(GIATRI_MOD)
	BEGIN
		CASE GIATRI_MOD IS
			WHEN "01" => DAU_CHAM_8LED <= X"FE";
			WHEN "10" => DAU_CHAM_8LED <= X"F7";
			WHEN OTHERS => DAU_CHAM_8LED <= X"FF";
		END CASE;
	END PROCESS;
		ENA_GIAIMA_8LED <= ENAGM_8LED_REG;
end Behavioral;

