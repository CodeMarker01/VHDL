library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity Bai8_3chuongtrinh is
	Port ( CKHT: in STD_LOGIC;
			BTN: IN STD_LOGIC_VECTOR(1 DOWNTO 0);
			LED: out STD_LOGIC_VECTOR (7 downto 0));
end Bai8_3chuongtrinh;

architecture Behavioral of Bai8_3chuongtrinh is
SIGNAL RST,ENA_DB,CHEDO: STD_LOGIC;
SIGNAL Q_STD,Q_SDTH_TSP,Q_4TRAI_4PHAI: STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL MODE: STD_LOGIC_VECTOR(2 DOWNTO 0);
Begin
	RST <= NOT BTN(0);
	CHEDO <= NOT BTN(1);
	
CHIA_10ENA: ENTITY WORK.CHIA_10ENA
	PORT MAP ( CKHT => CKHT,
	ENA5HZ => ENA_DB);
	
LED8_STD_PST: ENTITY WORK.LED8_STD_PST
	PORT MAP ( CKHT => CKHT,
	RST => RST,
	ENA_DB => ENA_DB,
	Q => Q_STD);
	

LED8_SDTH_TSP: ENTITY WORK.LED8_SDTH_TSP
	PORT MAP ( CKHT => CKHT,
	RST => RST,
	ENA_DB => ENA_DB,
	Q => Q_SDTH_TSP);
	
LED8_4TRAI_4PHAI: ENTITY WORK.LED8_4TRAI_4PHAI
	PORT MAP ( CKHT => CKHT,
	RST => RST,
	ENA_DB => ENA_DB,
	Q => Q_4TRAI_4PHAI);
	
DEM_3BIT_BTN: ENTITY WORK.DEM_3BIT_BTN
	PORT MAP ( CKHT => CKHT,
	RST => RST,
	BTN => CHEDO,
	Q => MODE);
	
LED <= Q_STD WHEN MODE ="001" ELSE
		 Q_4TRAI_4PHAI WHEN MODE ="010" ELSE
		 Q_SDTH_TSP WHEN MODE ="011" ELSE
		 "00000000";
		 
	
end Behavioral;