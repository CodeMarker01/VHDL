library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity DEM_4BIT_BTN is
	Port ( CKHT, RST, BTN: in STD_LOGIC;
			Q: out STD_LOGIC_VECTOR (3 downto 0));
end DEM_4BIT_BTN;

architecture Behavioral of DEM_4BIT_BTN is
SIGNAL ENA_DB: STD_LOGIC;
BEGIN
	CD_LAM_HEP_BTN: ENTITY WORK.CD_LAM_HEP_BTN
	PORT MAP ( CKHT => CKHT,
	BTN => BTN,
	BTN_CDLH => ENA_DB);
	DEM_4BIT: ENTITY WORK.DEM_4BIT
	PORT MAP ( CKHT => CKHT,
	RST => RST,
	ENA_DB => ENA_DB,
	Q => Q);
end Behavioral;