
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity DEM_4BIT_DK is
    Port (CKHT,RST, BTN_UP,BTN_DW,BTN_XUNG, ENA10HZ,ENA1HZ,ENA2HZ,ENA5HZ,ENA20HZ: in  STD_LOGIC;
				ENA_DB: OUT STD_LOGIC;
    		Q:    out    STD_LOGIC_VECTOR (3 downto 0));
end DEM_4BIT_DK;

architecture Behavioral of DEM_4BIT_DK is
SIGNAL 	Q_REG, Q_NEXT: STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL 	Q1_REG, Q1_NEXT: STD_LOGIC_VECTOR(3 DOWNTO 0);
BEGIN
	PROCESS (CKHT )
	BEGIN	
		
		IF	FALLING_EDGE (CKHT)  THEN  	Q_REG	<=	Q_NEXT;	
		END IF;
	END PROCESS;
	PROCESS (CKHT,RST )
	BEGIN	
		IF RST ='1' THEN  Q1_REG	<=	"0000";	
		ELSIF	FALLING_EDGE (CKHT)  THEN  	Q1_REG	<=	Q1_NEXT;	
		END IF;
	END PROCESS;
	
	Q_NEXT <= 	"0011" WHEN BTN_UP = '1'	AND Q_REG="1111" ELSE
					Q_REG+1 WHEN BTN_UP = '1' ELSE
					"1111" WHEN BTN_DW = '1'	AND Q_REG="0011" ELSE
					Q_REG -1 WHEN BTN_DW = '1'	 ELSE
					Q_REG ; 					
	Q	<= Q_REG;
	Q1_NEXT <= "0000"WHEN BTN_XUNG='1' AND Q1_REG ="0100" ELSE 
					Q1_REG+1 WHEN BTN_XUNG='1' ELSE
					Q1_REG;
	ENA_DB<= ENA1HZ WHEN Q1_REG ="0000" ELSE
				ENA2HZ WHEN Q1_REG ="0001" ELSE 
				ENA5HZ WHEN Q1_REG ="0010" ELSE 
				ENA10HZ WHEN Q1_REG ="0011" ELSE 
				ENA20HZ ;	
end Behavioral;

