LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY DEM_8BIT IS
	PORT(CKHT,RST, ENA_DB:IN STD_LOGIC;
			SS: OUT STD_LOGIC;
			PST_TSP: OUT STD_LOGIC_VECTOR(1 DOWNTO 0)
			);
END DEM_8BIT;

ARCHITECTURE BEHAVIORAL OF DEM_8BIT IS
SIGNAL Q_REG,Q_NEXT : STD_LOGIC_VECTOR(7 DOWNTO 0);
BEGIN
	PROCESS(CKHT,RST)
	BEGIN
		IF(RST='1') THEN Q_REG <= (OTHERS=>'0');
		ELSIF FALLING_EDGE(CKHT) THEN Q_REG <= Q_NEXT;
		END IF;
	END PROCESS;
	Q_NEXT <=  X"01" 			WHEN ENA_DB = '1' AND Q_REG =X"04" ELSE
				Q_REG+1     WHEN ENA_DB='1' 						  ELSE 
				 Q_REG;	
	SS<= '0' WHEN Q_REG =X"02" OR Q_REG =X"04" OR Q_REG=X"00" ELSE 
			'1';
	PST_TSP<= 	"01" WHEN Q_REG =X"01" OR Q_REG =X"02"ELSE 
					"10" WHEN Q_REG =X"03" OR Q_REG =X"04" ELSE 
					"00" ;
					
										
END BEHAVIORAL;