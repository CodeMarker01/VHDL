
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity GIA_TRI_CAI_NHAP_NHAY is
    Port ( CKHT : in  STD_LOGIC;
           BELL : out  STD_LOGIC;
           BTN_N : in  STD_LOGIC_VECTOR (4 downto 0);
           ANODE, SSEG : out  STD_LOGIC_VECTOR (7 downto 0));
end GIA_TRI_CAI_NHAP_NHAY;

architecture Behavioral of GIA_TRI_CAI_NHAP_NHAY is

SIGNAL ENA_DB, ENA1KHZ, ENA2HZ, ENA_CHINH, RST, BTN_DW, BTN_UP, BTN_SS, BTN_MOD : STD_LOGIC;

SIGNAL GIAY, PHUT, GIAY_CHINH, PHUT_CHINH: STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL CH_PHUT, DV_PHUT: STD_LOGIC_VECTOR (3 DOWNTO 0);
SIGNAL CH_GIAY, DV_GIAY: STD_LOGIC_VECTOR (3 DOWNTO 0);

SIGNAL CH_PHUT_CHINH, DV_PHUT_CHINH: STD_LOGIC_VECTOR (3 DOWNTO 0);
SIGNAL CH_GIAY_CHINH, DV_GIAY_CHINH: STD_LOGIC_VECTOR (3 DOWNTO 0);

SIGNAL LED0, LED1, LED2, LED3: STD_LOGIC_VECTOR (3 DOWNTO 0);


SIGNAL ENA_SS, ENA_DW, ENA_NN, ENA_UP: STD_LOGIC;

SIGNAL GIATRI_MOD: STD_LOGIC_VECTOR( 1 DOWNTO 0);
SIGNAL DAU_CHAM_8LED: STD_LOGIC_VECTOR (7 DOWNTO 0);
SIGNAL ENA_GIAIMA_8LED: STD_LOGIC_VECTOR (7 DOWNTO 0);
begin
	BELL <= '1';
	RST <= NOT BTN_N(0);
	BTN_DW <= NOT BTN_N(1);
	BTN_UP <= NOT BTN_N(2);
	BTN_MOD <= NOT BTN_N(3);
	BTN_SS <= NOT BTN_N(4);
	
CHIA_10ENA: ENTITY WORK.CHIA_10ENA
			PORT MAP(	CKHT => CKHT,
							ENA5HZ => ENA_DB,
							ENA10HZ => ENA2HZ,
							ENA1KHZ => ENA1KHZ);
							
CHONGDOI_DW: ENTITY WORK.DEBOUNCE_BTN
			PORT MAP(	CKHT => CKHT,
							BTN => BTN_DW,
							DB_TICK => ENA_DW);	
							
CHONGDOI_UP: ENTITY WORK.DEBOUNCE_BTN
			PORT MAP(	CKHT => CKHT,
							BTN => BTN_UP,
							DB_TICK => ENA_UP);	
							
NUT_NHAN_SS: ENTITY WORK.DEM_1BIT_BTN
			PORT MAP(	CKHT => CKHT,
							RST => RST,
							BTN => BTN_SS,
							Q => ENA_SS);
							
NUT_NHAN_MOD: ENTITY WORK.DEM_2BIT_BTN
			PORT MAP(	CKHT => CKHT,
							RST => RST,
							BTN => BTN_MOD,
							Q => GIATRI_MOD);
							
DEMXUONG_PHUTGIAY: ENTITY WORK.DEM_GIOPHUTGIAY
			PORT MAP(	CKHT => CKHT,
							RST => RST,
							ENA_NN => ENA_NN,
							ENA_DB => ENA_DB,
							ENA_SS => ENA_SS,
							ENA_UP => ENA_UP,
							ENA_DW => ENA_DW,
							ENA2HZ => ENA2HZ,
							GIATRI_MOD => GIATRI_MOD,
							PHUT => PHUT,
							GIAY => GIAY);
									
XULY_MOD_DAUCHAM_NHAP_NHAY:	ENTITY WORK.XULY_MOD_DAUCHAM_NHAP_NHAY
			PORT MAP(	CKHT => CKHT,
							ENA_DB => ENA_DB,
							ENA2HZ => ENA2HZ,
							ENA_DW => ENA_DW,
							ENA_UP => ENA_UP,
							ENA_NN => ENA_NN,
							ENA_SS => ENA_SS,
							ENA_GIAIMA_8LED => ENA_GIAIMA_8LED,
							GIATRI_MOD => GIATRI_MOD,
							DAU_CHAM_8LED => DAU_CHAM_8LED);
							

HEXTOBCD_PHUT: ENTITY WORK.HEXTOBCD_6BIT
			PORT MAP(	SOHEX6BIT => PHUT,
							DONVI => DV_PHUT,
							CHUC => CH_PHUT);
							
HEXTOBCD_GIAY: ENTITY WORK.HEXTOBCD_6BIT
			PORT MAP(	SOHEX6BIT => GIAY,
							DONVI => DV_GIAY,
							CHUC => CH_GIAY);
							
HIENTHI_2LED: ENTITY WORK.GIAIMA_HIENTHI_8LED_7DOAN
			PORT MAP(
					CKHT => CKHT,
					ENA1KHZ => ENA1KHZ,
					LED70 => DV_GIAY,
					LED71 => CH_GIAY, --- NHO SUA CHO NAY
					LED72 => X"F",
					LED73 => DV_PHUT,
					LED74 => CH_PHUT,
					LED75 => X"F",
					LED76 => X"F",
					LED77 => X"F",
					DAU_CHAM_8LED => DAU_CHAM_8LED,
					ENA_GIAIMA_8LED => ENA_GIAIMA_8LED,
					ANODE => ANODE,
					SSEG => SSEG);			
end Behavioral;

