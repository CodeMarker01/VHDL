LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY DEM_GIAY IS
	PORT(CKHT,RST, ENA_DB,ENA1HZ,ENA2HZ,ENA4HZ:IN STD_LOGIC;
			ENA_KQ: OUT STD_LOGIC);
END DEM_GIAY;

ARCHITECTURE BEHAVIORAL OF DEM_GIAY IS
SIGNAL Q_REG,Q_NEXT : STD_LOGIC_VECTOR(7 DOWNTO 0);
BEGIN
	PROCESS(CKHT,RST)
	BEGIN
		IF(RST='1') THEN Q_REG <= (OTHERS=>'0');
		ELSIF FALLING_EDGE(CKHT) THEN Q_REG <= Q_NEXT;
		END IF;
	END PROCESS;
	Q_NEXT <= Q_REG+1 WHEN ENA_DB ='1' AND Q_REG < 6 ELSE
				 Q_REG;
	--Q      <= Q_REG;
	ENA_KQ<= ENA1HZ WHEN Q_REG <2 ELSE
				ENA2HZ WHEN Q_REG <4 ELSE
				ENA4HZ;
END BEHAVIORAL;