-- CHUONG TRINH CON
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
entity MOD50_UD_CHILD is
Port ( CKHT, RST, ENA_DB, ENA_UD: in STD_LOGIC;
		 Q: out STD_LOGIC_VECTOR (5 downto 0);
		 SW: IN STD_LOGIC
		 );
end MOD50_UD_CHILD;
architecture Behavioral of MOD50_UD_CHILD is
SIGNAL Q_REG, Q_NEXT: STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL TEMP_Q_REG : STD_LOGIC_VECTOR (5 DOWNTO 0);
BEGIN
	PROCESS (CKHT, RST,SW)
		BEGIN
		-- NEU RESET = 1 THI GAN NGO RA = 0
			IF RST='1' AND SW='0' THEN Q_REG <= (OTHERS => '0'); --ENA_UD <= '0';
			ELSIF RST='1' AND SW='1' THEN Q_REG <= "110001"; --ENA_UD <= '1';
			ELSIF FALLING_EDGE (CKHT) THEN Q_REG <= Q_NEXT;
			ELSE 
		END IF;
	END PROCESS;
	-- MOD 50
	TEMP_Q_REG <= (OTHERS => '0') WHEN ENA_UD = '1' AND Q_REG = "110010" ELSE
					  "110001" WHEN ENA_UD = '0' AND Q_REG = "111111" ELSE
					  Q_REG + 1 WHEN ENA_UD = '0' OR SW = '0' ELSE
					  Q_REG - 1 WHEN ENA_UD = '1' OR SW = '1' ELSE
					  Q_REG;
--	-- SW
--	PROCESS (SW)
--	BEGIN
--		IF SW = '0' THEN ENA_UD <= '0';
--		ELSE 				  ENA_UD <= '1';
--		END IF;
--	END PROCESS;

	Q_NEXT <= TEMP_Q_REG WHEN ENA_DB = '1' ELSE
				 Q_REG;
	Q <= Q_REG;
end Behavioral;