LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY DEM_NHI_PHAN_8BIT_UD_4CD IS
	PORT(CKHT, BTN_N0,BTN_N1:IN STD_LOGIC;
				LEDR: OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END DEM_NHI_PHAN_8BIT_UD_4CD;

ARCHITECTURE BEHAVIORAL OF DEM_NHI_PHAN_8BIT_UD_4CD IS
SIGNAL ENA_DB,RST,CD,DK,UP_DOWN,SS,ENA1HZ,ENA5HZ : STD_LOGIC;
BEGIN
	RST <= NOT BTN_N0;
	CD <= NOT BTN_N1;
CHIA_10ENA: ENTITY WORK.CHIA_10ENA
		PORT MAP ( CKHT => CKHT,
						ENA1HZ=>ENA1HZ,
						ENA5HZ=>ENA5HZ);
CD_LAM_HEP_BTN: ENTITY WORK.CD_LAM_HEP_BTN
PORT MAP (
					CKHT => CKHT,
					BTN=>CD,
					BTN_CDLH=> DK
			);		
DEM_8BIT: ENTITY WORK.DEM_8BIT
		PORT MAP (CKHT => CKHT,
						RST => RST,
						ENA_DB=> DK,
						CK1HZ=>ENA1HZ,
						CK5HZ=>ENA5HZ,
						UP_DOWN=>UP_DOWN,
						SS => SS,
						ENA_KQ=>ENA_DB
					);			
DEM_8BIT_UD_SS: ENTITY WORK.DEM_8BIT_UD_SS
		PORT MAP (CKHT => CKHT,
						RST => RST,
						ENA_DB=> ENA_DB,
						ENA_SS=>SS,
						ENA_UD => UP_DOWN,
						Q => LEDR);
END BEHAVIORAL;