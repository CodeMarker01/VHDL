
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity DEM_0_15_0_10_0 is
		PORT(
					CKHT, BTN_N0: IN STD_LOGIC;
					BELL: OUT STD_LOGIC;
					ENA_SS: IN STD_LOGIC;
					LED_N: OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
			);
end DEM_0_15_0_10_0;

architecture Behavioral of DEM_0_15_0_10_0 is
SIGNAL ENA_DB, RST, ENA_UD, STATE: STD_LOGIC;
SIGNAL DK_STATE : STD_LOGIC_VECTOR(1 DOWNTO 0);
SIGNAL LED: STD_LOGIC_VECTOR(3 DOWNTO 0);
begin
		BELL <= '1';
		LED_N <= NOT LED; 
		RST <= NOT BTN_N0;

CHIA_10ENA: ENTITY WORK.CHIA_10ENA
	PORT MAP (
					CKHT => CKHT,
					ENA2HZ => ENA_DB
				);
				
DEM_4BIT: ENTITY WORK.DEM_8BIT  --4 BIT
	PORT MAP(
					CKHT => CKHT,
					RST => RST,
					ENA_DB => ENA_DB,
					ENA_UD => ENA_UD,
					ENA_SS => ENA_SS,
					STATE => STATE,
					Q => LED
				);	

STATE_DKHIEN: ENTITY WORK.STATE_DKHIEN
	PORT MAP(
					CKHT => CKHT,
					RST => RST,
					DK_STATE => DK_STATE,
					STATE => LED,
					Q_DKHIEN => ENA_UD					
				);	

DEM_2BIT: ENTITY WORK.DEM_2BIT
	PORT MAP(
					CKHT => CKHT,
					RST => RST,
					ENA_DB => ENA_DB,
					STATE => STATE,
					Q => DK_STATE					
				);	
 
end Behavioral;

