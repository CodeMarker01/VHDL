library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
entity HEXTOBCD_4BIT is
Port ( 	SOHEX4BIT: in STD_LOGIC_VECTOR (3 downto 0);
			DONVI, CHUC: out STD_LOGIC_VECTOR (3 downto 0));
end HEXTOBCD_4BIT;
architecture Behavioral of HEXTOBCD_4BIT is
BEGIN
	PROCESS (SOHEX4BIT)
	VARIABLE BCD_HEX: STD_LOGIC_VECTOR(11 DOWNTO 0);
	VARIABLE DEM: INTEGER RANGE 0 TO 3 ;
	BEGIN
		BCD_HEX:= "00000000" & SOHEX4BIT;
		DEM:= 3;
		WHILE DEM > 0
		LOOP
			BCD_HEX:= BCD_HEX(10 DOWNTO 0) & BCD_HEX(11);
			DEM:= DEM - 1;
			IF BCD_HEX(7 DOWNTO 4)>= "0101" THEN
				BCD_HEX(7 DOWNTO 4):= BCD_HEX(7 DOWNTO 4)+"0011";
			END IF;
			IF BCD_HEX(11 DOWNTO 8)>= "0101" THEN
				BCD_HEX(11 DOWNTO 8):= BCD_HEX(11 DOWNTO 8)+"0011";
			END IF;
		END LOOP;
		BCD_HEX:= BCD_HEX(10 DOWNTO 0) & '0';
		DONVI <= BCD_HEX(7 DOWNTO 4);
		CHUC <= BCD_HEX(11 DOWNTO 8);
	END PROCESS;
end Behavioral;