
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity LED8_4TRAI_4PHAI is
	Port ( CKHT, RST: in STD_LOGIC;
			ENA_DB: in STD_LOGIC;
			Q: out STD_LOGIC_VECTOR (7 downto 0));
end LED8_4TRAI_4PHAI;

architecture Behavioral of LED8_4TRAI_4PHAI is
SIGNAL Q_REG, Q_NEXT,Q_TAM: STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL DEM_REG, DEM_NEXT: INTEGER RANGE 0 TO 10:=0;
Begin
	PROCESS (CKHT, RST)
	BEGIN
		IF RST='1' THEN Q_REG <= (OTHERS => '0');
							 DEM_REG <=0;
		ELSIF FALLING_EDGE (CKHT) THEN Q_REG <= Q_NEXT;
												 DEM_REG <= DEM_NEXT;
		END IF;
	END PROCESS;
	
	DEM_NEXT <= 0 WHEN DEM_REG = 9 AND ENA_DB ='1' ELSE	
				DEM_REG + 1 WHEN ENA_DB ='1' ELSE
				DEM_REG;
				
	PROCESS (DEM_NEXT)
	BEGIN
				IF DEM_REG =0 THEN Q_NEXT <= (OTHERS => '1');
		ELSIF DEM_REG = 1 THEN Q_NEXT <= (OTHERS => '0');
		ELSIF DEM_REG = 2 THEN Q_NEXT <= (OTHERS => '1');
		ELSIF DEM_REG = 3 THEN Q_NEXT <= (OTHERS => '0');
		ELSIF DEM_REG = 4 THEN Q_NEXT <= (OTHERS => '1');
		ELSIF DEM_REG = 5 THEN Q_NEXT <= (OTHERS => '0');
		ELSIF DEM_REG = 6 THEN Q_NEXT <= "11110000";
		ELSIF DEM_REG = 7 THEN Q_NEXT <= (OTHERS => '0');
		ELSIF DEM_REG = 8 THEN Q_NEXT <= "11110000";
		ELSIF DEM_REG = 9 THEN Q_NEXT <= (OTHERS => '0');
		END IF;
	END PROCESS;
	
	
----------------------	

	Q <= Q_REG ;
end Behavioral;