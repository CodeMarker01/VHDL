
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity DEM_6BIT is
    Port ( CKHT : in  STD_LOGIC;
           ENA_DB : in  STD_LOGIC;
           ENA_SS1, ENA_SS2, ENA_SS3, ENA_SS4 : in  STD_LOGIC;
           Q : out  STD_LOGIC_VECTOR (5 downto 0));
end DEM_6BIT;

architecture Behavioral of DEM_6BIT is
signal Q_NEXT1: STD_LOGIC_VECTOR(5 DOWNTO 0);
signal Q_NEXT2: STD_LOGIC_VECTOR(5 DOWNTO 0);
signal Q_NEXT3: STD_LOGIC_VECTOR(5 DOWNTO 0);
signal Q_NEXT4: STD_LOGIC_VECTOR(5 DOWNTO 0);


signal Q_REG1: STD_LOGIC_VECTOR(5 DOWNTO 0):="000001";
signal Q_REG2: STD_LOGIC_VECTOR(5 DOWNTO 0):="000110";
signal Q_REG3: STD_LOGIC_VECTOR(5 DOWNTO 0):="001011";
signal Q_REG4: STD_LOGIC_VECTOR(5 DOWNTO 0):="010000";

begin
PROCESS(CKHT)
	BEGIN
		IF FALLING_EDGE (CKHT) THEN Q_REG1 <= Q_NEXT1;
											Q_REG2 <= Q_NEXT2;
											Q_REG3 <= Q_NEXT3;
											Q_REG4 <= Q_NEXT4;
		END IF;
	END PROCESS;
	
PROCESS(ENA_DB, ENA_SS1, ENA_SS2, ENA_SS3, ENA_SS4, Q_REG1, Q_REG2, Q_REG3, Q_REG4)	
	BEGIN
		IF (ENA_DB = '1' AND ENA_SS1 ='1' AND ENA_SS2 ='0' AND ENA_SS3 ='0' AND ENA_SS4='0') THEN
				Q_NEXT1 <= Q_REG1 +1;
			 IF Q_REG1 = "110011" THEN 
				Q_NEXT1 <="000001";
			END IF;
				Q <= Q_REG1;
		ELSIF (ENA_DB = '1' AND ENA_SS2 ='1' AND ENA_SS1 ='0' AND ENA_SS3 ='0' AND ENA_SS4='0') THEN
				Q_NEXT2 <= Q_REG2 + 1;
			 IF Q_REG2 = "110011" THEN 
				Q_NEXT2 <="000110" ;
			END IF;
				Q <= Q_REG2;
		ELSIF (ENA_DB = '1' AND ENA_SS3 ='1' AND ENA_SS2 ='0' AND ENA_SS1 ='0' AND ENA_SS4='0') THEN
				Q_NEXT3 <= Q_REG3 +1;
			 IF Q_REG3 = "110011" THEN 
				 Q_NEXT3 <="001011";
			END IF;
				Q <= Q_REG3;
		ELSIF (ENA_DB = '1' AND ENA_SS4 ='1' AND ENA_SS2 ='0' AND ENA_SS3 ='0' AND ENA_SS1='0') THEN
				Q_NEXT4 <= Q_REG4 +1;
			 IF Q_REG4 = "110011" THEN 
				Q_NEXT4 <="010000";
			END IF;
				Q <= Q_REG4;
		END IF;
	END PROCESS;
			
end Behavioral;