library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity DEM_8BIT_SS is
Port (CKHT, RST, ENA_DB,ENA_SS: in STD_LOGIC;
Q: out STD_LOGIC_VECTOR (7 downto 0));
end DEM_8BIT_SS;

architecture Behavioral of DEM_8BIT_SS is
SIGNAL Q_REG, Q_NEXT: STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL ENA_TMP:STD_LOGIC;
BEGIN
ENA_TMP <=ENA_DB;
	PROCESS (CKHT, RST)
	BEGIN
		IF ENA_SS='0' THEN ENA_TMP <= '0' ;
		ELSIF RST='1' THEN Q_REG <= (OTHERS => '0');
		ELSIF FALLING_EDGE (CKHT) THEN Q_REG <= Q_NEXT;
		END IF;
	END PROCESS;
	Q_NEXT <= Q_REG + 1 WHEN ENA_DB = '1' ELSE
	Q_REG;
	Q <= Q_REG;
end Behavioral;