library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity DIEUKHIEN_CHOPHEP is
Port ( CKHT, RST, ENA_DB: in STD_LOGIC;
OE: out STD_LOGIC_VECTOR (3 downto 0));
end DIEUKHIEN_CHOPHEP;

architecture Behavioral of DIEUKHIEN_CHOPHEP is
SIGNAL DEM_REG, DEM_NEXT: INTEGER RANGE 0 TO 47:=0;
begin
	PROCESS(CKHT, RST)
	BEGIN
		IF (RST ='1') THEN DEM_REG <= 0;
		ELSIF FALLING_EDGE(CKHT) THEN DEM_REG <= DEM_NEXT;
		END IF;
	END PROCESS;
	DEM_NEXT <= 0 WHEN DEM_REG = 47 AND ENA_DB = '1' ELSE
	DEM_REG + 1 WHEN ENA_DB = '1' ELSE
	DEM_REG;
	PROCESS(DEM_REG)
	BEGIN
		OE <= "0000";
		IF DEM_REG < 16 THEN OE <= "0001";
		ELSIF DEM_REG < 32 THEN OE <= "0010";
		ELSIF DEM_REG < 40 THEN OE <= "0100";
		ELSIF DEM_REG < 48 THEN OE <= "1000";
		END IF;
	END PROCESS;
end Behavioral;