-- TAO XUNG TICH CUC MUC 1 DUNG BANG 1 CHU KI ckth
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
entity CHIA_1ENA1HZ is
	Port ( CKHT: in STD_LOGIC;
			ENA1HZ: out STD_LOGIC);
end CHIA_1ENA1HZ;
architecture Behavioral of CHIA_1ENA1HZ is
CONSTANT N: INTEGER:= 50000000;
SIGNAL D1HZ_REG, D1HZ_NEXT: INTEGER RANGE 0 TO N:=1;
Begin
	PROCESS (CKHT)
	BEGIN
	-- REGISTER: NEU CO XUNG THI GAN
		IF FALLING_EDGE (CKHT) THEN D1HZ_REG <= D1HZ_NEXT;
		END IF;
	END PROCESS;
	-- D1HZ_REG = N THI GAN D1HZ_NEXT = 1 -> CHU KI MOI
	-- NEU KO THI D1HZ_REG + 1
	D1HZ_NEXT <= 1 WHEN D1HZ_REG = N ELSE
					 D1HZ_REG + 1;
	-- ENA1HZ CHI BANG 1 KHI D1HZ_REG DUNG = N/2
	ENA1HZ <= '1' WHEN D1HZ_REG = N/2 ELSE '0';
end Behavioral;