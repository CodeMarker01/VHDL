library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity DEM_8BIT_SS_UD_AUTO is
Port (CKHT, RST, ENA_DB,ENA_SS: in STD_LOGIC;
Q: out STD_LOGIC_VECTOR (7 downto 0));
end DEM_8BIT_SS_UD_AUTO;

architecture Behavioral of DEM_8BIT_SS_UD_AUTO is
SIGNAL Q_REG, Q_NEXT_UP,Q_NEXT_DW,Q_TMP: STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL ENA_TMP,TMP:STD_LOGIC;

BEGIN
ENA_TMP <=ENA_DB;
	PROCESS (CKHT, RST)
	BEGIN
		IF ENA_SS='0' THEN ENA_TMP <= '0' ;
		ELSIF RST='1' THEN Q_REG <= (OTHERS => '0');
		ELSIF FALLING_EDGE (CKHT) THEN Q_REG <= Q_TMP;
		END IF;
	END PROCESS;
	
	PROCESS (Q_REG)
	BEGIN
		IF Q_REG="11111111" THEN TMP <='0';
		ELSIF Q_REG="00000000" THEN TMP <='1';
		END IF;
	END PROCESS;
	
	Q_TMP <= Q_NEXT_UP WHEN TMP='1' ELSE	
				Q_NEXT_DW;
	
	Q_NEXT_UP <= Q_REG + 1 WHEN ENA_DB = '1'  ELSE
	Q_REG;
	
	Q_NEXT_DW <= Q_REG - 1 WHEN ENA_DB = '1'  ELSE
	Q_REG;
	
	Q <= Q_REG;
end Behavioral;