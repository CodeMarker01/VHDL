-- CHUONG TRINH CON
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;

entity CHIA_2XUNG is
Port ( CKHT: in STD_LOGIC;
		CK1HZ,CK10HZ: out STD_LOGIC);
end CHIA_2XUNG;

architecture Behavioral of CHIA_2XUNG is
CONSTANT N: INTEGER := 50000000;
-- 1 XUNG CK -> 1 HZ
SIGNAL D1HZ_REG, D1HZ_NEXT: INTEGER RANGE 0 TO N:=1;
-- 10 XUNG CK -> 1 HZ
SIGNAL D10HZ_REG, D10HZ_NEXT: INTEGER RANGE 0 TO N/10:=1;
Begin
	--REGISTER D-FF
	PROCESS (CKHT)
	BEGIN
		IF FALLING_EDGE (CKHT) THEN D1HZ_REG <= D1HZ_NEXT;
											 D10HZ_REG <= D10HZ_NEXT;
		END IF;
	END PROCESS;
		--NEXT STATE LOGIC
		D1HZ_NEXT <= 1 WHEN D1HZ_REG = N ELSE
						 D1HZ_REG + 1;
		D10HZ_NEXT <= 1 WHEN D1HZ_REG = N/10 ELSE
						 D10HZ_REG +1;
		
		--OUTOUT LOGIC
		CK1HZ <= '1' WHEN D1HZ_REG < N/2 ELSE
					'0';
		CK10HZ <= '1' WHEN D1HZ_REG < N/20 ELSE
					 '0';
end Behavioral;