-- DEM LEN 8 BIT
-- RESET MUC 1
-- ENA_SS MUC 1: DEM, MUC 0: NGUNG
-- ENA_UD : 1 LEN, 0 XUONG
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
entity DEM_MOD40_UD is
Port ( CKHT: in STD_LOGIC;
		LED: out STD_LOGIC_VECTOR (5 downto 0);
		SW: in STD_LOGIC_VECTOR(1 DOWnto 0);
		BTN_N: IN STD_LOGIC_VECTOR(1 DOWnto 0));
end DEM_MOD40_UD;
architecture Behavioral of DEM_MOD40_UD is
SIGNAL ENA_DB, RST: STD_LOGIC;
SIGNAL ENA_UD: STD_LOGIC;
begin
	RST <= NOT BTN_N(0);
--	ENA_UD <= NOT BTN_N(1);
--	CHIA_1ENA1HZ: ENTITY WORK.CHIA_10ENA
	CHIA_1ENA1HZ: ENTITY WORK.CHIA_10ENA
	PORT MAP ( CKHT => CKHT,
				  ena5hz => ENA_DB);
	DEM_1BIT_BTN: ENTITY WORK.DEM_1BIT
	PORT MAP ( CKHT => CKHT,
					RST => RST,
				  ENA_DB => ENA_DB,
				  Q => ENA_UD);
	CD_LAM_HEP_BTN: ENTITY WORK.CD_LAM_HEP_BTN
	PORT MAP ( CKHT => CKHT,
					BTN => BTN_N(1),
					BTN_CDLH => ENA_DB);
	DEM_8BIT: ENTITY WORK.DEM_MOD40_UD_CTC
	PORT MAP ( CKHT => CKHT,
					RST => RST,
					ENA_DB => ENA_DB,
					Q => LED,
					ENA_SS => SW(0),
					ENA_UD => ENA_UD);
end Behavioral;