library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity DEM_6BIT is
	Port ( CKHT: in STD_LOGIC;
			 ENA_DB_UP, ENA_DB_DW: in STD_LOGIC;
			 UP, DW: IN STD_LOGIC;
			 ENA_UP, ENA_DW: IN STD_LOGIC;
			Q: out STD_LOGIC_VECTOR (5 downto 0));
end DEM_6BIT;

architecture Behavioral of DEM_6BIT is
SIGNAL Q_REG, Q_NEXT: STD_LOGIC_VECTOR(5 DOWNTO 0);
BEGIN
	PROCESS (CKHT, UP, DW)
	BEGIN
--		IF RST='1' THEN Q_REG <= (OTHERS => '0');
		IF UP = '1' THEN Q_REG <= "000001";
		ELSIF DW = '1' THEN Q_REG <= "111111";
		ELSIF FALLING_EDGE (CKHT) THEN Q_REG <= Q_NEXT;
		END IF;
	END PROCESS;
	Q_NEXT <= Q_REG + 1 WHEN ENA_DB_UP = '1' AND ENA_UP = '1' ELSE
				 Q_REG - 1 WHEN ENA_DB_DW = '1' AND ENA_DW = '1' ELSE
				 Q_REG;
	Q <= Q_REG;
end Behavioral;