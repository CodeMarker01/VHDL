library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity DIEUKHIEN_CHOPHEP is
	Port ( CKHT, RST, ENA_DB: in STD_LOGIC;
			OE: out STD_LOGIC_VECTOR (7 downto 0));
end DIEUKHIEN_CHOPHEP;

architecture Behavioral of DIEUKHIEN_CHOPHEP is
SIGNAL DEM_REG, DEM_NEXT: INTEGER RANGE 0 TO 137:=0;
begin
	PROCESS(CKHT, RST)
	BEGIN
		IF (RST ='1') THEN DEM_REG <= 0;
		ELSIF FALLING_EDGE(CKHT) THEN DEM_REG <= DEM_NEXT;
		END IF;
	END PROCESS;
	DEM_NEXT <= 0 WHEN DEM_REG = 137 AND ENA_DB = '1' ELSE
	DEM_REG + 1 WHEN ENA_DB = '1' ELSE
	DEM_REG;
	PROCESS(DEM_REG)
	BEGIN
	
		OE <= "00000000";
		IF DEM_REG < 16 THEN OE <= "00000001";
		ELSIF DEM_REG < 32 THEN OE <= "00000010";
		ELSIF DEM_REG < 40 THEN OE <= "00000100";
		ELSIF DEM_REG < 48 THEN OE <= "00001000";
		ELSIF DEM_REG < 56 THEN OE <= "00010000";
		ELSIF DEM_REG < 64 THEN OE <= "00100000";
		ELSIF DEM_REG < 101 THEN OE <= "01000000";
		ELSIF DEM_REG < 138 THEN OE <= "10000000";
		END IF;
		
	END PROCESS;
end Behavioral;