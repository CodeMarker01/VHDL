library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
entity DK_8LED_SELECT_STD_PST_TSP is
Port ( CKHT,BTN_N0,SW0: in STD_LOGIC;
LED: out STD_LOGIC_VECTOR (7 downto 0));
end DK_8LED_SELECT_STD_PST_TSP;
architecture Behavioral of DK_8LED_SELECT_STD_PST_TSP is
SIGNAL ENA_DB, RST: STD_LOGIC;
SIGNAL Q_STD_PST, Q_STD_TSP: STD_LOGIC_VECTOR (7 downto 0);
SIGNAL OE: STD_LOGIC_VECTOR(1 DOWNTO 0);
Begin
RST <= NOT BTN_N0;
CHIA_10ENA: ENTITY WORK.CHIA_10ENA
	PORT MAP ( CKHT => CKHT,
					ENA5HZ => ENA_DB);
LED_STD_PST: ENTITY WORK.LED_STD_PST
	PORT MAP ( CKHT => CKHT,
					RST => RST,
					ENA_DB => ENA_DB,
					OE => OE(0),
					Q => Q_STD_PST);
LED_STD_TSP: ENTITY WORK.LED_STD_TSP
	PORT MAP ( CKHT => CKHT,
					RST => RST,
					ENA_DB => ENA_DB,
					OE => OE(1),
					Q => Q_STD_TSP);
LED <= Q_STD_PST OR Q_STD_TSP;
OE <= "01" WHEN SW0='0' ELSE
"10";
end Behavioral;