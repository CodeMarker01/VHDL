
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;



entity THAY_DOI_TAN_SO is
    Port ( CKHT, BTN_N0 : in  STD_LOGIC;
           BELL : out  STD_LOGIC;
           ANODE, SSEG : out  STD_LOGIC_VECTOR (7 downto 0));
end THAY_DOI_TAN_SO;

architecture Behavioral of THAY_DOI_TAN_SO is
SIGNAL ENA_DB, ENA1HZ, ENA2HZ, ENA5HZ, ENA10HZ, ENA1KHZ, RST: STD_LOGIC;
SIGNAL DONVI, CHUC: STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL S: STD_LOGIC_VECTOR(1 DOWNTO 0);
SIGNAL DEM: STD_LOGIC_VECTOR(5 DOWNTO 0):="000001";
SIGNAL DAU_CHAM_8LED: STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL ENA_GIAIMA_8LED: STD_LOGIC_VECTOR(7 DOWNTO 0);

begin

	BELL <= '1';
	RST <= NOT BTN_N0;
	DAU_CHAM_8LED <= X"FF";
	ENA_GIAIMA_8LED <= X"07";	
	
CHIA_10ENA: ENTITY WORK.CHIA_10ENA
			PORT MAP(	CKHT => CKHT,
							ENA1HZ => ENA1HZ,
							ENA5HZ => ENA2HZ,
							ENA10HZ => ENA5HZ,
							ENA20HZ => ENA10HZ,
							ENA1KHZ => ENA1KHZ);	
							
CHON_TAN_SO: ENTITY WORK.CHON_TAN_SO
			PORT MAP(	CKHT => CKHT,
							RST => RST,
							CHUC => CHUC,
							DONVI => DONVI,
							Q => S);
							
	ENA_DB  <=  ENA1HZ WHEN S = "00" ELSE
					ENA2HZ WHEN S = "01" ELSE
					ENA5HZ WHEN S = "10" ELSE
					ENA10HZ;	
					
DEM_0_50: ENTITY WORK.DEM_6BIT
			PORT MAP(	CKHT => CKHT,
							RST => RST,
							ENA_DB => ENA_DB,
							Q => DEM);
							
HEXTOBCD: ENTITY WORK.HEXTOBCD_6BIT
			PORT MAP(	SOHEX6BIT => DEM,
							DONVI => DONVI,
							CHUC => CHUC);
							
HIENTHI_2LED: ENTITY WORK.GIAIMA_HIENTHI_8LED_7DOAN
			PORT MAP(
					CKHT => CKHT,
					ENA1KHZ => ENA1KHZ,
					LED70 => DONVI,
					LED71 => CHUC,
					LED72 => X"F",
					LED73 => X"F",
					LED74 => X"F",
					LED75 => X"F",
					LED76 => X"F",
					LED77 => X"F",
					DAU_CHAM_8LED => DAU_CHAM_8LED,
					ENA_GIAIMA_8LED => ENA_GIAIMA_8LED,
					ANODE => ANODE,
					SSEG => SSEG);
end Behavioral;

