
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity GIO_NHIET_DO is
    Port ( CKHT : in  STD_LOGIC;
           BELL : out  STD_LOGIC;
           BTN_N : in  STD_LOGIC_VECTOR (1 downto 0);
           DS18B20 : inout  STD_LOGIC;
			  DECIMAL : out  STD_LOGIC_VECTOR (3 downto 0);
           SSEG, ANODE : out  STD_LOGIC_VECTOR (7 downto 0));
end GIO_NHIET_DO;

architecture Behavioral of GIO_NHIET_DO is
SIGNAL ENA_DB, ENA1KHZ, RST, BTN_MOD, Q, DS_PRESENT : STD_LOGIC;
SIGNAL GIAY, PHUT, GIO: STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL GIO5: STD_LOGIC_VECTOR (4 DOWNTO 0);

SIGNAL CH_GIO, DV_GIO: STD_LOGIC_VECTOR (3 DOWNTO 0);
SIGNAL CH_PHUT, DV_PHUT: STD_LOGIC_VECTOR (3 DOWNTO 0);
SIGNAL CH_GIAY, DV_GIAY: STD_LOGIC_VECTOR (3 DOWNTO 0);

SIGNAL DAU_CHAM_8LED: STD_LOGIC_VECTOR (7 DOWNTO 0);
SIGNAL ENA_GIAIMA_8LED: STD_LOGIC_VECTOR (7 DOWNTO 0);

SIGNAL DONVI, CHUC, TRAM: STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL LED0, LED1, LED2: STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL LED_0, LED_1, LED_2, LED_3, LED_4, LED_5, LED_6, LED_7: STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL NHIETDO: STD_LOGIC_VECTOR (7 DOWNTO 0);
SIGNAL TEMPERATURE: STD_LOGIC_VECTOR (11 DOWNTO 0);

begin

	RST <= NOT BTN_N(0);
	BTN_MOD <= NOT BTN_N(1);
	DAU_CHAM_8LED <= X"FF";
	ENA_GIAIMA_8LED <= "11011011" WHEN Q ='1' ELSE "11000111";
	GIO <= '0'& GIO5;
	BELL <= '0' WHEN (DONVI >= 2 AND CHUC >= 3) ELSE '1';
CHIA_10ENA: ENTITY WORK.CHIA_10ENA
			PORT MAP(	CKHT => CKHT,
							ENA20HZ => ENA_DB,
							ENA1KHZ => ENA1KHZ);
							
NUT_MOD: ENTITY WORK.DEM_1BIT_BTN
			PORT MAP(	CKHT => CKHT,
							RST => RST,
							BTN => BTN_MOD,
							Q => Q);
							
DEM_GIOPHUTGIAY: ENTITY WORK.DEM_GIOPHUTGIAY
			PORT MAP(	CKHT => CKHT,
							RST => RST,
							ENA_DB => ENA_DB,
							GIO => GIO5,
							PHUT => PHUT,
							GIAY => GIAY);
HEXTOBCD_GIO: ENTITY WORK.HEXTOBCD_6BIT
			PORT MAP(	SOHEX6BIT => GIO,
							DONVI => DV_GIO,
							CHUC => CH_GIO);
							
HEXTOBCD_PHUT: ENTITY WORK.HEXTOBCD_6BIT
			PORT MAP(	SOHEX6BIT => PHUT,
							DONVI => DV_PHUT,
							CHUC => CH_PHUT);
							
HEXTOBCD_GIAY: ENTITY WORK.HEXTOBCD_6BIT
			PORT MAP(	SOHEX6BIT => GIAY,
							DONVI => DV_GIAY,
							CHUC => CH_GIAY);
---------------------------------------------------------------------------
NHIETDO <= TEMPERATURE (11 DOWNTO 4);
DECIMAL <= TEMPERATURE (3 DOWNTO 0);
	
DS18B20_TEMPERATURE: ENTITY WORK.DS18B20_TEMPERATURE
	PORT MAP ( 	CKHT => CKHT,
					RST => RST,
					DS18B20 => DS18B20,
					DS_PRESENT => DS_PRESENT,
					TEMPERATURE_OUT => TEMPERATURE);
	PROCESS (DS_PRESENT, DONVI, CHUC, TRAM)
	BEGIN
		IF (DS_PRESENT = '0') THEN
									LED0 <= DONVI;
									LED1 <= CHUC;
									LED2 <= TRAM;
		ELSE
									LED0 <= X"E";
									LED1 <= X"E";
									LED2 <= X"E";
		END IF;
	END PROCESS;
	
	
						
HEXTOBCD_ND: ENTITY WORK.HEXTOBCD_8BIT
			PORT MAP(	SOHEX8BIT => NHIETDO,
							DONVI => DONVI,
							CHUC => CHUC,
							TRAM => TRAM);		
---------------------------------------------------------------------------	
LED_0 <= DV_GIAY WHEN Q = '1' ELSE LED0;
LED_1 <= CH_GIAY WHEN Q = '1' ELSE LED1;
LED_2 <= X"F" WHEN Q = '1' ELSE LED2;
LED_3 <= DV_PHUT WHEN Q = '1' ELSE X"F";
LED_4 <= CH_PHUT WHEN Q = '1' ELSE X"F";
LED_5 <= X"F" WHEN Q = '1' ELSE X"F";
LED_6 <= DV_GIO WHEN Q = '1' ELSE X"2";
LED_7 <= CH_GIO WHEN Q = '1' ELSE X"3";
---------------------------------------------------------------------------					
HIENTHI_2LED: ENTITY WORK.GIAIMA_HIENTHI_8LED_7DOAN
			PORT MAP(
					CKHT => CKHT,
					ENA1KHZ => ENA1KHZ,
					LED70 => LED_0,
					LED71 => LED_1, --- NHO SUA CHO NAY
					LED72 => LED_2,
					LED73 => LED_3,
					LED74 => LED_4,
					LED75 => LED_5,
					LED76 => LED_6,
					LED77 => LED_7,
					DAU_CHAM_8LED => DAU_CHAM_8LED,
					ENA_GIAIMA_8LED => ENA_GIAIMA_8LED,
					ANODE => ANODE,
					SSEG => SSEG);										

end Behavioral;

