LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY DEM_8BIT IS
	PORT(CKHT,RST, ENA_DB:IN STD_LOGIC;
			SW: IN STD_LOGIC_VECTOR(2 DOWNTO 0);
			SO_LED: OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
			);
END DEM_8BIT;

ARCHITECTURE BEHAVIORAL OF DEM_8BIT IS
SIGNAL Q_REG,Q_NEXT : STD_LOGIC_VECTOR(7 DOWNTO 0);
BEGIN
	PROCESS(CKHT,RST)
	BEGIN
		IF(RST='1') 					THEN Q_REG <= (OTHERS=>'0');
		ELSIF FALLING_EDGE(CKHT)   THEN Q_REG <= Q_NEXT;
		END IF;
	END PROCESS;
	Q_NEXT <=  X"00" WHEN ENA_DB ='1' AND Q_REG=X"03"  ELSE
				  X"01" WHEN ENA_DB ='1' AND SW="000" 		ELSE
				  X"02" WHEN ENA_DB ='1' AND SW="001"  	ELSE					 
				  X"03" WHEN ENA_DB ='1' AND SW="011" 		ELSE
				  Q_REG;
				 
	SO_LED<= "0011" WHEN Q_REG=X"01" AND  SW="001" ELSE
				"0111" WHEN Q_REG=X"02" AND  SW="011" ELSE
				"1111" WHEN Q_REG=X"03" AND  SW="111" ELSE
				"0001";
	--Q      <= Q_REG;
END BEHAVIORAL;