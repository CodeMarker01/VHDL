---- CHUONG TRINH CON
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
entity DEM_BIN_0_20_UP is
Port ( CKHT, RST, ENA_DB: in STD_LOGIC;
		 --OE: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		 OE: IN STD_LOGIC;
		 Q: out STD_LOGIC_VECTOR (5 downto 0));
end DEM_BIN_0_20_UP;
architecture Behavioral of DEM_BIN_0_20_UP is
SIGNAL Q_REG, Q_NEXT: STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL TEMP_Q_REG : STD_LOGIC_VECTOR (5 DOWNTO 0);
BEGIN
	PROCESS (CKHT, RST)
		BEGIN
		-- NEU RESET = 1 THI GAN NGO RA = 0
			IF RST='1' THEN Q_REG <= (OTHERS => '0');
			ELSIF FALLING_EDGE (CKHT) THEN Q_REG <= Q_NEXT;
			ELSE 
		END IF;
	END PROCESS;
	Q_NEXT <= (OTHERS => '0') WHEN Q_REG = "101001" ELSE
					  Q_REG + 1 WHEN ENA_DB = '1' AND OE = '1' ELSE
					  Q_REG;
	Q <= Q_REG;
end Behavioral;