library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;

entity CHIA_1ENA1HZ is
Port ( CKHT: in STD_LOGIC;
		ENA1HZ: out STD_LOGIC);
end CHIA_1ENA1HZ;

architecture Behavioral of CHIA_1ENA1HZ is
CONSTANT N: INTEGER:= 50000000;
SIGNAL D1HZ_REG, D1HZ_NEXT: INTEGER RANGE 0 TO N:=1;
Begin
	PROCESS (CKHT)
	BEGIN
	-- D-FF: CO XUNG THI GAN
		IF FALLING_EDGE (CKHT) THEN D1HZ_REG <= D1HZ_NEXT;
		END IF;
	END PROCESS;
	-- HET 50M XUNG THI RESET VE 1
	-- CHUA HET 50M XUNG THI TIEP TUC CONG
	D1HZ_NEXT <= 1 WHEN D1HZ_REG = N ELSE
					 D1HZ_REG + 1;
	-- TAI DUNG N/2 THI LEN MUC 1 (CUC NHANH)
	ENA1HZ <= '1' WHEN D1HZ_REG = N/2 ELSE '0';
end Behavioral;