
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;


entity XULY_MOD_DAUCHAM_NHAP_NHAY is
    Port ( CKHT, ENA_DB, ENA2HZ, ENA_UP, ENA_DW, ENA_HT, RST, SS_ND : in  STD_LOGIC;
           GIATRI_MOD : out  STD_LOGIC_VECTOR (1 downto 0);
           ENA_GIAIMA_8LED,NHIET_DO, GIOI_HAN_ND : out  STD_LOGIC_VECTOR (7 downto 0);
           DAU_CHAM_8LED : out  STD_LOGIC_VECTOR (7 downto 0));
end XULY_MOD_DAUCHAM_NHAP_NHAY;

architecture Behavioral of XULY_MOD_DAUCHAM_NHAP_NHAY is
SIGNAL GIATRI_MOD_REG: STD_LOGIC_VECTOR( 1 DOWNTO 0):="00";
SIGNAL GIATRI_MOD_NEXT: STD_LOGIC_VECTOR( 1 DOWNTO 0);
SIGNAL ENAGM_8LED_REG: STD_LOGIC_VECTOR( 7 DOWNTO 0):=X"FF";
SIGNAL ENAGM_8LED_NEXT: STD_LOGIC_VECTOR( 7 DOWNTO 0);
SIGNAL DLNN_REG: STD_LOGIC_VECTOR( 4 DOWNTO 0):="00000";
SIGNAL DLNN_NEXT: STD_LOGIC_VECTOR( 4 DOWNTO 0);

begin
	PROCESS(CKHT)
	BEGIN
		IF FALLING_EDGE(CKHT) THEN GIATRI_MOD_REG <= GIATRI_MOD_NEXT;
											ENAGM_8LED_REG <= ENAGM_8LED_NEXT;
											DLNN_REG <= DLNN_NEXT;
		END IF;
	END PROCESS;
	GIATRI_MOD_NEXT <= GIATRI_MOD_REG + 1 WHEN (ENA_DB = '1' AND ENA_HT ='0') ELSE
								"00" WHEN (DLNN_REG = "10100" OR RST ='1' OR ENA_HT ='1') ELSE --CHO NAY LA KHI DLNN = 20 THI SE K EDIT DC TIME LED SE K NN NUA
								GIATRI_MOD_REG;
	PROCESS(GIATRI_MOD_REG, ENA_UP, ENA_DW, ENA2HZ, ENAGM_8LED_REG, DLNN_REG, ENA_HT, SS_ND)
	BEGIN
		ENAGM_8LED_NEXT <= ENAGM_8LED_REG;
		DLNN_NEXT <= DLNN_REG;
		IF GIATRI_MOD_REG = "01" AND ENA_HT = '0' THEN
			IF (ENA_UP = '0' AND ENA_DW = '0') THEN
				IF ENA2HZ = '1' THEN 
					ENAGM_8LED_NEXT <= "110110" & NOT ENAGM_8LED_REG( 1 DOWNTO 0); --NHAP NHAY 2 LED GIAY
					DLNN_NEXT <= DLNN_REG + 1; --DEM THOI GIAN NHAP NHAY
				END IF;
			ELSE
				ENAGM_8LED_NEXT <= X"DB"; --CAC LED SANG BT 11011011
				DLNN_NEXT <= (OTHERS => '0'); --NEU UP OR DW = 1 THI RESET BIEN DEM NN
			END IF;
		
		-----------------------------------------------------------------------
		ELSIF GIATRI_MOD_REG = "10" AND ENA_HT = '0' THEN
			IF (ENA_UP = '0' AND ENA_DW = '0') THEN
				IF ENA2HZ = '1' THEN 
					ENAGM_8LED_NEXT <= "110" & NOT ENAGM_8LED_REG( 4 DOWNTO 3) & "011"; --NHAP NHAY 2 LED PHUT
					DLNN_NEXT <= DLNN_REG + 1; --DEM THOI GIAN NHAP NHAY
				END IF;
			ELSE
				ENAGM_8LED_NEXT <= X"DB"; --CAC LED SANG BT 11011011
				DLNN_NEXT <= (OTHERS => '0'); --NEU UP OR DW = 1 THI RESET BIEN DEM NN
			END IF;
		----------------------------------------------------------------------------------------------
		ELSIF GIATRI_MOD_REG = "11" AND ENA_HT = '0' THEN
			IF (ENA_UP = '0' AND ENA_DW = '0') THEN
				IF ENA2HZ = '1' THEN 
					ENAGM_8LED_NEXT <= NOT ENAGM_8LED_REG( 7 DOWNTO 6) & "011011"; --NHAP NHAY 2 LED GIO
					DLNN_NEXT <= DLNN_REG + 1; --DEM THOI GIAN NHAP NHAY
				END IF;
			ELSE
				ENAGM_8LED_NEXT <= X"DB"; --CAC LED SANG BT 11011011
				DLNN_NEXT <= (OTHERS => '0'); --NEU UP OR DW = 1 THI RESET BIEN DEM NN
			END IF;
		----------------------------------------------------------------------------------------------
		ELSIF GIATRI_MOD_REG = "00" AND ENA_HT = '1' THEN
			IF SS_ND = '1' THEN
				IF ENA2HZ = '1' THEN 
					ENAGM_8LED_NEXT <= NOT ENAGM_8LED_REG( 7 DOWNTO 6) & "0000" & NOT ENAGM_8LED_REG( 1 DOWNTO 0);
				END IF;
			ELSE
				ENAGM_8LED_NEXT <= "11000011";
			END IF;
		ELSE
				ENAGM_8LED_NEXT <= X"DB"; --CAC LED SANG BT 11011011
				DLNN_NEXT <= (OTHERS => '0'); --NEU UP OR DW = 1 THI RESET BIEN DEM NN
		END IF;
	END PROCESS;
		
		------------------------------------------------------------
		
		DAU_CHAM_8LED <= X"FE" WHEN GIATRI_MOD_REG = "01" AND ENA_HT ='0' ELSE
							  X"F7" WHEN GIATRI_MOD_REG = "10" AND ENA_HT ='0' ELSE
							  X"BF" WHEN GIATRI_MOD_REG = "11" AND ENA_HT ='0' ELSE
							  X"FF";
							  
		GIATRI_MOD <= GIATRI_MOD_REG;
		ENA_GIAIMA_8LED <= ENAGM_8LED_REG;
end Behavioral;

