
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;


entity TOI_GOIHAN_XX is
    Port ( CKHT, SW0 : in  STD_LOGIC;
           BTN_N : in  STD_LOGIC_VECTOR (1 downto 0);
           SSEG, ANODE : out  STD_LOGIC_VECTOR (7 downto 0);
           BELL : out  STD_LOGIC);
end TOI_GOIHAN_XX;

architecture Behavioral of TOI_GOIHAN_XX is

SIGNAL ENA_DB, ENA1KHZ, RST, BTN: STD_LOGIC;
SIGNAL DONVI, CHUC, TRAM, DONVI_XX, CHUC_XX, TRAM_XX: STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL DEM: STD_LOGIC_VECTOR(7 DOWNTO 0):=X"00";
SIGNAL DAU_CHAM_8LED: STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL GH: STD_LOGIC_VECTOR(7 DOWNTO 0);

SIGNAL Q: STD_LOGIC_VECTOR(1 DOWNTO 0);
SIGNAL ENA_GIAIMA_8LED: STD_LOGIC_VECTOR(7 DOWNTO 0);

begin
	BELL <= '1';
	RST <= NOT BTN_N(0);
	BTN <= NOT BTN_N(1);
	DAU_CHAM_8LED <= X"FF";
	
XOA_SO_0: ENTITY WORK.XOA_SO_0_VN
			PORT MAP(	CHUC => CHUC,
							TRAM => TRAM,
							ENA_GIAIMA_8LED => ENA_GIAIMA_8LED);
							
CHIA_10ENA: ENTITY WORK.CHIA_10ENA
			PORT MAP(	CKHT => CKHT,
							ENA2HZ => ENA_DB,
							ENA1KHZ => ENA1KHZ);	
							
NUT_NHAN_GH: ENTITY WORK.DEM_2BIT_BTN
			PORT MAP(	CKHT => CKHT,
							RST => RST,
							BTN => BTN,
							Q => Q);
 GH <= "01011010" WHEN Q ="00"	ELSE
			"01010000" WHEN Q ="01" ELSE
			"01000110" WHEN Q ="10" ELSE
			"00111100";						
			
DEM_200_XX: ENTITY WORK.DEM_8BIT
			PORT MAP(	CKHT => CKHT,
							RST => RST,
							ENA_DB => ENA_DB,
							GH => GH,
							DEM => DEM);
							
HEXTOBCD: ENTITY WORK.HEXTOBCD_8BIT
			PORT MAP(	SOHEX8BIT => DEM,
							DONVI => DONVI,
							CHUC => CHUC,
							TRAM => TRAM);
HEXTOBCD_HT: ENTITY WORK.HEXTOBCD_8BIT
			PORT MAP(	SOHEX8BIT => GH,
							DONVI => DONVI_XX,
							CHUC => CHUC_XX,
							TRAM => TRAM_XX);
							
HIENTHI_2LED: ENTITY WORK.GIAIMA_HIENTHI_8LED_7DOAN
			PORT MAP(
					CKHT => CKHT,
					ENA1KHZ => ENA1KHZ,
					LED70 => DONVI,
					LED71 => CHUC, --- NHO SUA CHO NAY
					LED72 => TRAM,
					LED73 => X"F",
					LED74 => X"F",
					LED75 => X"F",
					LED76 => DONVI_XX,
					LED77 => CHUC_XX,
					DAU_CHAM_8LED => DAU_CHAM_8LED,
					ENA_GIAIMA_8LED => ENA_GIAIMA_8LED,
					ANODE => ANODE,
					SSEG => SSEG);

end Behavioral;

