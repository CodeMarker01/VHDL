LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY DEM_8BIT IS
	PORT(CKHT,RST, ENA_DB:IN STD_LOGIC;
			Q: OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END DEM_8BIT;

ARCHITECTURE BEHAVIORAL OF DEM_8BIT IS
SIGNAL Q_REG,Q_NEXT : STD_LOGIC_VECTOR(7 DOWNTO 0);
BEGIN
	PROCESS(CKHT,RST)
	BEGIN
		IF(RST='1') THEN Q_REG <= (OTHERS=>'0');
		ELSIF FALLING_EDGE(CKHT) THEN Q_REG <= Q_NEXT;
		END IF;
	END PROCESS;
	Q_NEXT <= Q_REG+1 WHEN ENA_DB ='1' ELSE
				 Q_REG;
	Q      <= Q_REG;
END BEHAVIORAL;