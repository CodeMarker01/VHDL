-- CHUONG TRINH CON
-- ENA_DB : 
-- ENA_SS : CHO PHEP DEM HAY NGUNG DEM
-- ENA_UD : CHO PHEP DEM LEN HAY DEM XUONG
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
entity DEM_8BIT_SS_UD_AUTO is
-- BO ENA_UD
Port ( CKHT, RST, ENA_DB, ENA_SS: in STD_LOGIC;
		 Q: out STD_LOGIC_VECTOR (7 downto 0));
end DEM_8BIT_SS_UD_AUTO;
architecture Behavioral of DEM_8BIT_SS_UD_AUTO is
SIGNAL Q_REG, Q_NEXT: STD_LOGIC_VECTOR(7 DOWNTO 0);
--SIGNAL TEMP_Q_REG : STD_LOGIC_VECTOR (7 DOWNTO 0);
--SIGNAL TEMP_COUNT : STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL ENA_UD_REG, ENA_UD_NEXT: STD_LOGIC;
BEGIN
	PROCESS (CKHT, RST)
		BEGIN
		-- NEU RESET = 1 THI GAN NGO RA = 0
			IF RST='1' THEN Q_REG <= (OTHERS => '0');
								 ENA_UD_REG <= '0'; -- MACH DEM LEN KHI NHAN RESET
			ELSIF FALLING_EDGE (CKHT) THEN Q_REG <= Q_NEXT;
											ENA_UD_REG <= ENA_UD_NEXT;
		END IF;
	END PROCESS;
--	ENA_UD_NEXT <= '1' WHEN Q_REG = "11111111" ELSE
--						'0' WHEN Q_REG = "00000000" ELSE
--						ENA_UD_REG;
	
--	TEMP_Q_REG <= Q_REG + 1 WHEN ENA_UD_REG = '0' ELSE
--					  Q_REG - 1;

	Q_NEXT <= Q_REG + 1 WHEN ENA_DB = '1' AND ENA_SS='1' AND ENA_UD_REG = '0' ELSE
				 Q_REG - 1 WHEN ENA_DB = '1' AND ENA_SS='1' AND ENA_UD_REG = '1' ELSE
				 Q_REG;
	Q <= Q_REG;
end Behavioral;